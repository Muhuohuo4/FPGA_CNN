module conv11_input #(
    parameter DATA_WIDTH = 8
)(
    input  wire clk,
    input  wire rst,

    // 来自滑窗的数据输入
    input  wire input_valid,
    input  wire inputbuf_read_en,
    input  wire [DATA_WIDTH-1:0] data_in,

    // 输出给卷积计算模块
    output wire [DATA_WIDTH-1:0] out_0_0,

    // 控制信号输出
    output wire input_ready
);

    // 中间信号
    wire inputbuf_load;

    // 数据缓存模块实例化
    conv11_input_buffer #(
        .DATA_WIDTH(DATA_WIDTH)
    ) u_input_buffer (
        .clk(clk),
        .rst(rst),
        .input_valid(input_valid),
        .inputbuf_read_en(inputbuf_read_en),
        .inputbuf_load(inputbuf_load),
        .data_in(data_in),
        .out_0_0(out_0_0)
    );

    // 控制模块实例化
    conv11_input_ctrl u_input_ctrl (
        .clk(clk),
        .rst(rst),
        .input_valid(input_valid),
        .inputbuf_load(inputbuf_load),
        .input_ready(input_ready)
    );

endmodule
