module channel_2 #(parameter DEPTH = 16900) (
    input  wire        clk,
    input  wire        we,
    input  wire [13:0] addr_write,
    input  wire [13:0] addr_read,
    input  wire [7:0]  data_in,
    output wire [7:0]  data_out
);
    (* ram_style = "block" *) reg [7:0] mem [0:DEPTH-1];
    initial $readmemh("G.mem", mem);  // 仿真用
    
    always @(posedge clk) begin
        if (we)
            mem[addr_write] <= data_in;
    end

    assign data_out = mem[addr_read];

endmodule
