module conv33_output_buffer #(
    parameter OUT_WIDTH = 32
)(
    input wire clk,
    input wire rst,

    // 来自计算模块的输出
    input wire in_valid,
    input wire [OUT_WIDTH-1:0] in_data, 

    // 控制模块指示何时读取
    input wire read_en,

    // 输出给下一模块
    output reg out_valid, 
    output reg [OUT_WIDTH-1:0] out_data 
);

    // 内部缓冲  
    reg [OUT_WIDTH-1:0] buffer;
    reg buffer_valid;

    // 写入缓冲
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            buffer <= 0;
            buffer_valid <= 0;
        end else if (in_valid) begin
            buffer <= in_data;
            buffer_valid <= 1;
        end else if (read_en) begin
            buffer_valid <= 0; 
        end
    end

    // 输出逻辑
    always @(posedge clk) begin
        if (read_en && buffer_valid) begin
            out_data  <= buffer;
            out_valid <= 1;
        end else begin
            out_valid <= 0;
        end
    end

endmodule
