module sliding_window_3x3 (
    input  wire        clk,
    input  wire        rst,
    input  wire        en,                    // 输入使能，每拍一个像素
    input  wire signed [7:0]  pixel_in,       // 输入像素
    output reg         valid,                 // 输出有效
    output reg  signed [7:0]  o_temp [0:8]    // 3x3 窗口：左上→右下
);

    parameter IMG_WIDTH = 130;

    // === 两行缓冲 ===
    reg signed [7:0] line_buf_0 [0:IMG_WIDTH-1];  // 行 n-2
    reg signed [7:0] line_buf_1 [0:IMG_WIDTH-1];  // 行 n-1

    reg signed [7:0] shift_col_0 [0:2];
    reg signed [7:0] shift_col_1 [0:2];
    reg signed [7:0] shift_col_2 [0:2];

    reg [13:0] col_cnt;
    reg [13:0] pix_cnt;

    // 计数器更新
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            col_cnt <= 0;
            pix_cnt <= 0;
        end else if (en) begin
            pix_cnt <= pix_cnt + 1;
            col_cnt <= (col_cnt == IMG_WIDTH-1) ? 0 : col_cnt + 1;
        end
    end

    // 行缓冲写入
    always @(posedge clk) begin
        if (en) begin
            line_buf_0[col_cnt] <= line_buf_1[col_cnt];
            line_buf_1[col_cnt] <= pixel_in;
        end
    end

    // 列移位
    always @(posedge clk) begin
        if (en) begin
            shift_col_0[0] <= shift_col_0[1];
            shift_col_0[1] <= shift_col_0[2];
            shift_col_0[2] <= line_buf_0 [col_cnt];

            shift_col_1[0] <= shift_col_1[1];
            shift_col_1[1] <= shift_col_1[2];
            shift_col_1[2] <= line_buf_1 [col_cnt];

            shift_col_2[0] <= shift_col_2[1];
            shift_col_2[1] <= shift_col_2[2];
            shift_col_2[2] <= pixel_in;
        end
    end

    // 拼窗口
    always @(posedge clk) begin
        if (en) begin
            o_temp[0] <= shift_col_0[0]; o_temp[1] <= shift_col_1[0]; o_temp[2] <= shift_col_2[0];
            o_temp[3] <= shift_col_0[1]; o_temp[4] <= shift_col_1[1]; o_temp[5] <= shift_col_2[1];
            o_temp[6] <= shift_col_0[2]; o_temp[7] <= shift_col_1[2]; o_temp[8] <= shift_col_2[2];
        end
    end

    // 有效信号
    always @(posedge clk or posedge rst) begin
        if (rst) valid <= 0;
        else     valid <= (en && pix_cnt >= IMG_WIDTH * 2 + 2);
    end


endmodule
