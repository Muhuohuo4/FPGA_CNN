`define CONV_0_IN_CHANNELS           3
`define CONV_0_OUT_CHANNELS          16
`define CONV_0_KERNEL_H              3
`define CONV_0_KERNEL_W              3
`define CONV_0_OUT_H                 64
`define CONV_0_OUT_W                 64
`define CONV_0_OUT_C                 16
`define CONV_0_STRIDE                1

`define CONV_DW_1_IN_CHANNELS        16
`define CONV_DW_1_OUT_CHANNELS       16
`define CONV_DW_1_KERNEL_H           3
`define CONV_DW_1_KERNEL_W           3
`define CONV_DW_1_OUT_H              64
`define CONV_DW_1_OUT_W              64
`define CONV_DW_1_OUT_C              16
`define CONV_DW_1_STRIDE             1

`define CONV_PW_1_IN_CHANNELS        16
`define CONV_PW_1_OUT_CHANNELS       32
`define CONV_PW_1_KERNEL_H           1
`define CONV_PW_1_KERNEL_W           1
`define CONV_PW_1_OUT_H              64
`define CONV_PW_1_OUT_W              64
`define CONV_PW_1_OUT_C              32
`define CONV_PW_1_STRIDE             1

`define CONV_DW_2_IN_CHANNELS        32
`define CONV_DW_2_OUT_CHANNELS       32
`define CONV_DW_2_KERNEL_H           3
`define CONV_DW_2_KERNEL_W           3
`define CONV_DW_2_OUT_H              32
`define CONV_DW_2_OUT_W              32
`define CONV_DW_2_OUT_C              32
`define CONV_DW_2_STRIDE             2

`define CONV_PW_2_IN_CHANNELS        32
`define CONV_PW_2_OUT_CHANNELS       64
`define CONV_PW_2_KERNEL_H           1
`define CONV_PW_2_KERNEL_W           1
`define CONV_PW_2_OUT_H              32
`define CONV_PW_2_OUT_W              32
`define CONV_PW_2_OUT_C              64
`define CONV_PW_2_STRIDE             1

`define CONV_DW_3_IN_CHANNELS        64
`define CONV_DW_3_OUT_CHANNELS       64
`define CONV_DW_3_KERNEL_H           3
`define CONV_DW_3_KERNEL_W           3
`define CONV_DW_3_OUT_H              32
`define CONV_DW_3_OUT_W              32
`define CONV_DW_3_OUT_C              64
`define CONV_DW_3_STRIDE             1

`define CONV_PW_3_IN_CHANNELS        64
`define CONV_PW_3_OUT_CHANNELS       64
`define CONV_PW_3_KERNEL_H           1
`define CONV_PW_3_KERNEL_W           1
`define CONV_PW_3_OUT_H              32
`define CONV_PW_3_OUT_W              32
`define CONV_PW_3_OUT_C              64
`define CONV_PW_3_STRIDE             1

`define CONV_DW_4_IN_CHANNELS        64
`define CONV_DW_4_OUT_CHANNELS       64
`define CONV_DW_4_KERNEL_H           3
`define CONV_DW_4_KERNEL_W           3
`define CONV_DW_4_OUT_H              16
`define CONV_DW_4_OUT_W              16
`define CONV_DW_4_OUT_C              64
`define CONV_DW_4_STRIDE             2

`define CONV_PW_4_IN_CHANNELS        64
`define CONV_PW_4_OUT_CHANNELS       128
`define CONV_PW_4_KERNEL_H           1
`define CONV_PW_4_KERNEL_W           1
`define CONV_PW_4_OUT_H              16
`define CONV_PW_4_OUT_W              16
`define CONV_PW_4_OUT_C              128
`define CONV_PW_4_STRIDE             1

`define CONV_DW_5_IN_CHANNELS        128
`define CONV_DW_5_OUT_CHANNELS       128
`define CONV_DW_5_KERNEL_H           3
`define CONV_DW_5_KERNEL_W           3
`define CONV_DW_5_OUT_H              16
`define CONV_DW_5_OUT_W              16
`define CONV_DW_5_OUT_C              128
`define CONV_DW_5_STRIDE             1

`define CONV_PW_5_IN_CHANNELS        128
`define CONV_PW_5_OUT_CHANNELS       128
`define CONV_PW_5_KERNEL_H           1
`define CONV_PW_5_KERNEL_W           1
`define CONV_PW_5_OUT_H              16
`define CONV_PW_5_OUT_W              16
`define CONV_PW_5_OUT_C              128
`define CONV_PW_5_STRIDE             1

`define CONV_DW_6_IN_CHANNELS        128
`define CONV_DW_6_OUT_CHANNELS       128
`define CONV_DW_6_KERNEL_H           3
`define CONV_DW_6_KERNEL_W           3
`define CONV_DW_6_OUT_H              16
`define CONV_DW_6_OUT_W              16
`define CONV_DW_6_OUT_C              128
`define CONV_DW_6_STRIDE             1

`define CONV_PW_6_IN_CHANNELS        128
`define CONV_PW_6_OUT_CHANNELS       128
`define CONV_PW_6_KERNEL_H           1
`define CONV_PW_6_KERNEL_W           1
`define CONV_PW_6_OUT_H              16
`define CONV_PW_6_OUT_W              16
`define CONV_PW_6_OUT_C              128
`define CONV_PW_6_STRIDE             1

`define CONV_DW_7_IN_CHANNELS        128
`define CONV_DW_7_OUT_CHANNELS       128
`define CONV_DW_7_KERNEL_H           3
`define CONV_DW_7_KERNEL_W           3
`define CONV_DW_7_OUT_H              16
`define CONV_DW_7_OUT_W              16
`define CONV_DW_7_OUT_C              128
`define CONV_DW_7_STRIDE             1

`define CONV_PW_7_IN_CHANNELS        128
`define CONV_PW_7_OUT_CHANNELS       128
`define CONV_PW_7_KERNEL_H           1
`define CONV_PW_7_KERNEL_W           1
`define CONV_PW_7_OUT_H              16
`define CONV_PW_7_OUT_W              16
`define CONV_PW_7_OUT_C              128
`define CONV_PW_7_STRIDE             1

`define CONV_DW_8_IN_CHANNELS        128
`define CONV_DW_8_OUT_CHANNELS       128
`define CONV_DW_8_KERNEL_H           3
`define CONV_DW_8_KERNEL_W           3
`define CONV_DW_8_OUT_H              16
`define CONV_DW_8_OUT_W              16
`define CONV_DW_8_OUT_C              128
`define CONV_DW_8_STRIDE             1

`define CONV_PW_8_IN_CHANNELS        128
`define CONV_PW_8_OUT_CHANNELS       128
`define CONV_PW_8_KERNEL_H           1
`define CONV_PW_8_KERNEL_W           1
`define CONV_PW_8_OUT_H              16
`define CONV_PW_8_OUT_W              16
`define CONV_PW_8_OUT_C              128
`define CONV_PW_8_STRIDE             1

`define CONV_DW_9_IN_CHANNELS        128
`define CONV_DW_9_OUT_CHANNELS       128
`define CONV_DW_9_KERNEL_H           3
`define CONV_DW_9_KERNEL_W           3
`define CONV_DW_9_OUT_H              16
`define CONV_DW_9_OUT_W              16
`define CONV_DW_9_OUT_C              128
`define CONV_DW_9_STRIDE             1

`define CONV_PW_9_IN_CHANNELS        128
`define CONV_PW_9_OUT_CHANNELS       128
`define CONV_PW_9_KERNEL_H           1
`define CONV_PW_9_KERNEL_W           1
`define CONV_PW_9_OUT_H              16
`define CONV_PW_9_OUT_W              16
`define CONV_PW_9_OUT_C              128
`define CONV_PW_9_STRIDE             1

`define CONV_DW_10_IN_CHANNELS       128
`define CONV_DW_10_OUT_CHANNELS      128
`define CONV_DW_10_KERNEL_H          3
`define CONV_DW_10_KERNEL_W          3
`define CONV_DW_10_OUT_H             8
`define CONV_DW_10_OUT_W             8
`define CONV_DW_10_OUT_C             128
`define CONV_DW_10_STRIDE            2

`define CONV_PW_10_IN_CHANNELS       128
`define CONV_PW_10_OUT_CHANNELS      256
`define CONV_PW_10_KERNEL_H          1
`define CONV_PW_10_KERNEL_W          1
`define CONV_PW_10_OUT_H             8
`define CONV_PW_10_OUT_W             8
`define CONV_PW_10_OUT_C             256
`define CONV_PW_10_STRIDE            1

`define CONV_DW_11_IN_CHANNELS       256
`define CONV_DW_11_OUT_CHANNELS      256
`define CONV_DW_11_KERNEL_H          3
`define CONV_DW_11_KERNEL_W          3
`define CONV_DW_11_OUT_H             8
`define CONV_DW_11_OUT_W             8
`define CONV_DW_11_OUT_C             256
`define CONV_DW_11_STRIDE            1

`define CONV_PW_11_IN_CHANNELS       256
`define CONV_PW_11_OUT_CHANNELS      256
`define CONV_PW_11_KERNEL_H          1
`define CONV_PW_11_KERNEL_W          1
`define CONV_PW_11_OUT_H             8
`define CONV_PW_11_OUT_W             8
`define CONV_PW_11_OUT_C             256
`define CONV_PW_11_STRIDE            1

`define CONV_DW_12_IN_CHANNELS       256
`define CONV_DW_12_OUT_CHANNELS      256
`define CONV_DW_12_KERNEL_H          3
`define CONV_DW_12_KERNEL_W          3
`define CONV_DW_12_OUT_H             4
`define CONV_DW_12_OUT_W             4
`define CONV_DW_12_OUT_C             256
`define CONV_DW_12_STRIDE            2

`define CONV_PW_12_IN_CHANNELS       256
`define CONV_PW_12_OUT_CHANNELS      512
`define CONV_PW_12_KERNEL_H          1
`define CONV_PW_12_KERNEL_W          1
`define CONV_PW_12_OUT_H             4
`define CONV_PW_12_OUT_W             4
`define CONV_PW_12_OUT_C             512
`define CONV_PW_12_STRIDE            1
