module conv11_bias_input #(
    parameter BIAS_WIDTH = 32
)(
    input  wire                  clk,
    input  wire                  rst,

    // 加载接口
    input  wire                  load_en,
    input  wire [BIAS_WIDTH-1:0] load_data,

    // 读取控制
    input  wire                  read_en,

    // 输出接口
    output reg  [BIAS_WIDTH-1:0] bias,        // 偏置输出
    output reg                   valid,       // 输出有效
    output reg                   bias_load    // 偏置加载完成（1拍脉冲）
);

    reg [BIAS_WIDTH-1:0] buffer;

    // 偏置加载过程
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            buffer     <= 0;
            bias_load  <= 0;
        end else if (load_en) begin
            buffer     <= load_data;
            bias_load  <= 1;  // 一拍脉冲，通知加载完成
        end else begin
            bias_load  <= 0;
        end
    end

    // 偏置读取输出
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            bias  <= 0;
            valid <= 0;
        end else if (read_en) begin
            bias  <= buffer;
            valid <= 1;
        end else begin
            valid <= 0;
        end
    end

endmodule
